`default_nettype none

module second ();
endmodule
